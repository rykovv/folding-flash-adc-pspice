** Profile: "SCHEMATIC1-testac"  [ C:\DOCUMENTS AND SETTINGS\PHEEDLEY\MY DOCUMENTS\PSPICE\EXAMPLES\EEE232\interp1\interp1-pspicefiles\schematic1\testac.sim ] 

** Creating circuit file "testac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../interp1-pspicefiles/interp1.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.01\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1k 10G
.OP
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
