** Profile: "SCHEMATIC1-testtran"  [ D:\OneDrive\OneDrive - Asian Answers\Documentos\CSUS\EEE232\Projects\Project 2\adc_flash_4b_interp_fold\adc_flash_4b_interp_fold-pspicefiles\schematic1\testtran.sim ] 

** Creating circuit file "testtran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../adc_flash_4b_interp_fold-pspicefiles/adc_flash_4b_interp_fold.lib" 
* From [PSPICE NETLIST] section of D:\Users\Vladmachine\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN/OP  0 10000n 0 0.5ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
